`include "uvm_macros.svh"  // Import UVM macros
import uvm_pkg::*;         // Import all UVM classes

parameter FIFO_DATA_WIDTH = 8;
`timescale 1ns / 1ps

/*
 * Acts as the FIFO Wrapper, that encapsulates all the FIFO components into a singular module that interacts with
 * the rx and tx mac via AXI Stream.
*/

module fifo
(

);
endmodule

`timescale 1ns / 1ps

module udp#(
    parameter AXI_DATA_WIDTH = 8
)(
    input wire i_clk,
    input wire i_reset_n,

    
);


endmodule : udp